library verilog;
use verilog.vl_types.all;
entity conv_tb is
end conv_tb;
