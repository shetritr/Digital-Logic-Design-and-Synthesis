library verilog;
use verilog.vl_types.all;
entity one_image_tb is
end one_image_tb;
