library verilog;
use verilog.vl_types.all;
entity TextFileReader_TB is
end TextFileReader_TB;
