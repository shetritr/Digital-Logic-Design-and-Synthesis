library verilog;
use verilog.vl_types.all;
entity CatRecognizer_tb is
end CatRecognizer_tb;
