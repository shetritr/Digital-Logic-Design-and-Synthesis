library verilog;
use verilog.vl_types.all;
entity Allimages_tb is
end Allimages_tb;
